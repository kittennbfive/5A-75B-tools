module top(input btn, output led);
	always begin
		led<=btn;
	end
endmodule
